module top();
      avalon_timer_qsys_tb tb ();
      test_program pgm ();
endmodule
