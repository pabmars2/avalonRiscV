// avalon_timer_qsys.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module avalon_timer_qsys (
		output wire  avalon_timer_0_external_interface_conduit, // avalon_timer_0_external_interface.conduit
		input  wire  clk_clk,                                   //                               clk.clk
		input  wire  reset_reset_n                              //                             reset.reset_n
	);

	wire  [31:0] mm_master_bfm_0_m0_readdata;                              // mm_interconnect_0:mm_master_bfm_0_m0_readdata -> mm_master_bfm_0:avm_readdata
	wire         mm_master_bfm_0_m0_waitrequest;                           // mm_interconnect_0:mm_master_bfm_0_m0_waitrequest -> mm_master_bfm_0:avm_waitrequest
	wire   [2:0] mm_master_bfm_0_m0_address;                               // mm_master_bfm_0:avm_address -> mm_interconnect_0:mm_master_bfm_0_m0_address
	wire         mm_master_bfm_0_m0_read;                                  // mm_master_bfm_0:avm_read -> mm_interconnect_0:mm_master_bfm_0_m0_read
	wire  [31:0] mm_master_bfm_0_m0_writedata;                             // mm_master_bfm_0:avm_writedata -> mm_interconnect_0:mm_master_bfm_0_m0_writedata
	wire         mm_master_bfm_0_m0_write;                                 // mm_master_bfm_0:avm_write -> mm_interconnect_0:mm_master_bfm_0_m0_write
	wire         mm_interconnect_0_avalon_timer_0_avalon_slave_chipselect; // mm_interconnect_0:avalon_timer_0_avalon_slave_chipselect -> avalon_timer_0:chipselect
	wire  [31:0] mm_interconnect_0_avalon_timer_0_avalon_slave_readdata;   // avalon_timer_0:readdata -> mm_interconnect_0:avalon_timer_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_avalon_timer_0_avalon_slave_address;    // mm_interconnect_0:avalon_timer_0_avalon_slave_address -> avalon_timer_0:address
	wire         mm_interconnect_0_avalon_timer_0_avalon_slave_read;       // mm_interconnect_0:avalon_timer_0_avalon_slave_read -> avalon_timer_0:read
	wire         mm_interconnect_0_avalon_timer_0_avalon_slave_write;      // mm_interconnect_0:avalon_timer_0_avalon_slave_write -> avalon_timer_0:write
	wire  [31:0] mm_interconnect_0_avalon_timer_0_avalon_slave_writedata;  // mm_interconnect_0:avalon_timer_0_avalon_slave_writedata -> avalon_timer_0:writedata
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> avalon_timer_0:reset
	wire         rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> [mm_interconnect_0:avalon_timer_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset, mm_master_bfm_0:reset]

	avalon_timer avalon_timer_0 (
		.clock      (clk_clk),                                                  //         clock_sink.clk
		.reset      (rst_controller_reset_out_reset),                           //         reset_sink.reset
		.irq        (),                                                         //   interrupt_sender.irq
		.chipselect (mm_interconnect_0_avalon_timer_0_avalon_slave_chipselect), //       avalon_slave.chipselect
		.address    (mm_interconnect_0_avalon_timer_0_avalon_slave_address),    //                   .address
		.write      (mm_interconnect_0_avalon_timer_0_avalon_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_avalon_timer_0_avalon_slave_writedata),  //                   .writedata
		.read       (mm_interconnect_0_avalon_timer_0_avalon_slave_read),       //                   .read
		.readdata   (mm_interconnect_0_avalon_timer_0_avalon_slave_readdata),   //                   .readdata
		.out_th     (avalon_timer_0_external_interface_conduit)                 // external_interface.conduit
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (3),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_master_bfm_0 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.avm_address            (mm_master_bfm_0_m0_address),         //        m0.address
		.avm_readdata           (mm_master_bfm_0_m0_readdata),        //          .readdata
		.avm_writedata          (mm_master_bfm_0_m0_writedata),       //          .writedata
		.avm_waitrequest        (mm_master_bfm_0_m0_waitrequest),     //          .waitrequest
		.avm_write              (mm_master_bfm_0_m0_write),           //          .write
		.avm_read               (mm_master_bfm_0_m0_read),            //          .read
		.avm_burstcount         (),                                   // (terminated)
		.avm_begintransfer      (),                                   // (terminated)
		.avm_beginbursttransfer (),                                   // (terminated)
		.avm_byteenable         (),                                   // (terminated)
		.avm_readdatavalid      (1'b0),                               // (terminated)
		.avm_arbiterlock        (),                                   // (terminated)
		.avm_lock               (),                                   // (terminated)
		.avm_debugaccess        (),                                   // (terminated)
		.avm_transactionid      (),                                   // (terminated)
		.avm_readid             (8'b00000000),                        // (terminated)
		.avm_writeid            (8'b00000000),                        // (terminated)
		.avm_clken              (),                                   // (terminated)
		.avm_response           (2'b00),                              // (terminated)
		.avm_writeresponsevalid (1'b0),                               // (terminated)
		.avm_readresponse       (8'b00000000),                        // (terminated)
		.avm_writeresponse      (8'b00000000)                         // (terminated)
	);

	avalon_timer_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                  //                                       clk_0_clk.clk
		.avalon_timer_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // avalon_timer_0_reset_sink_reset_bridge_in_reset.reset
		.mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // mm_master_bfm_0_clk_reset_reset_bridge_in_reset.reset
		.mm_master_bfm_0_m0_address                            (mm_master_bfm_0_m0_address),                               //                              mm_master_bfm_0_m0.address
		.mm_master_bfm_0_m0_waitrequest                        (mm_master_bfm_0_m0_waitrequest),                           //                                                .waitrequest
		.mm_master_bfm_0_m0_read                               (mm_master_bfm_0_m0_read),                                  //                                                .read
		.mm_master_bfm_0_m0_readdata                           (mm_master_bfm_0_m0_readdata),                              //                                                .readdata
		.mm_master_bfm_0_m0_write                              (mm_master_bfm_0_m0_write),                                 //                                                .write
		.mm_master_bfm_0_m0_writedata                          (mm_master_bfm_0_m0_writedata),                             //                                                .writedata
		.avalon_timer_0_avalon_slave_address                   (mm_interconnect_0_avalon_timer_0_avalon_slave_address),    //                     avalon_timer_0_avalon_slave.address
		.avalon_timer_0_avalon_slave_write                     (mm_interconnect_0_avalon_timer_0_avalon_slave_write),      //                                                .write
		.avalon_timer_0_avalon_slave_read                      (mm_interconnect_0_avalon_timer_0_avalon_slave_read),       //                                                .read
		.avalon_timer_0_avalon_slave_readdata                  (mm_interconnect_0_avalon_timer_0_avalon_slave_readdata),   //                                                .readdata
		.avalon_timer_0_avalon_slave_writedata                 (mm_interconnect_0_avalon_timer_0_avalon_slave_writedata),  //                                                .writedata
		.avalon_timer_0_avalon_slave_chipselect                (mm_interconnect_0_avalon_timer_0_avalon_slave_chipselect)  //                                                .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
