
module AvalonRiscV_QSYS (
	clk_clk,
	masteruart_rs232_rx_rx,
	masteruart_rs232_tx_tx,
	reset_reset_n);	

	input		clk_clk;
	input		masteruart_rs232_rx_rx;
	output		masteruart_rs232_tx_tx;
	input		reset_reset_n;
endmodule
