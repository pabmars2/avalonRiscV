
module avalon_timer_qsys (
	clk_clk,
	reset_reset_n,
	avalon_timer_0_external_interface_conduit);	

	input		clk_clk;
	input		reset_reset_n;
	output		avalon_timer_0_external_interface_conduit;
endmodule
