
module AvalonUARTQsys (
	avalon_timer_0_external_interface_conduit,
	avalonmasteruart_0_control_flag_tx,
	clk_clk,
	reset_reset_n);	

	output		avalon_timer_0_external_interface_conduit;
	input		avalonmasteruart_0_control_flag_tx;
	input		clk_clk;
	input		reset_reset_n;
endmodule
