module top();
      avalon_displays7seg_qsys_tb tb ();
      test_program pgm ();
endmodule
